module alu32_test;
    reg [31:0] A = 0, B = 0;
    reg [2:0] control = 0;

    initial begin
        $dumpfile("alu32.vcd");
        $dumpvars(0, alu32_test);

             A = 8; B = 4; control = `ALU_ADD; // try adding 8 and 4
        # 10 A = 2; B = 5; control = `ALU_SUB; // try subtracting 5 from 2

        # 10 A = 3; B = 4; control = `ALU_AND;
        # 10 A = 1; B = 5; control = `ALU_OR;
        # 10 A = 2; B = 3; control = `ALU_NOR;
        # 10 A = 6; B = 8; control = `ALU_XOR;

        # 10 A = 4; B = 4; control = `ALU_SUB;
        # 10 A = 32'h7ffffff0; B = 36; control = `ALU_SUB;


        # 10 A = 32'h7ffffff0; B = 32'h7fffffff; control = `ALU_ADD;
        # 10 A = 32'haffffff0; B = 32'hafffffff; control = `ALU_ADD;
        # 10 A = 32'h0ffffff0; B = 32'hfffffff0; control = `ALU_SUB;

        # 10 $finish;
    end

    wire [31:0] out;
    wire overflow, zero, negative;
    alu32 a(out, overflow, zero, negative, A, B, control);
endmodule // alu32_test
