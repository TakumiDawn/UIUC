// mips_decode: a decoder for MIPS arithmetic instructions
//
// alu_op       (output) - control signal to be sent to the ALU
// rd_src       (output) - should the destination register be rd (0) or rt (1)
// alu_src2     (output) - should the 2nd ALU source be a register (0) or an immediate (1)
// writeenable  (output) - should a new value be captured by the register file
// except       (output) - set to 1 when we don't recognize an opdcode & funct combination
// control_type (output) - 00 = fallthrough, 01 = branch_target, 10 = jump_target, 11 = jump_register
// mem_read     (output) - the register value written is coming from the memory
// word_we      (output) - we're writing a word's worth of data
// byte_we      (output) - we're only writing a byte's worth of data
// byte_load    (output) - we're doing a byte load
// slt          (output) - the instruction is an slt
// lui          (output) - the instruction is a lui
// addm         (output) - the instruction is an addm
// opcode        (input) - the opcode field from the instruction
// funct         (input) - the function field from the instruction
// zero          (input) - from the ALU
//

module mips_decode(alu_op, rd_src, alu_src2, writeenable, except, control_type,
                   mem_read, word_we, byte_we, byte_load, slt, lui, addm,
                   opcode, funct, zero);
    output [2:0] alu_op;
    output       rd_src, alu_src2, writeenable, except;
    output [1:0] control_type;
    output       mem_read, word_we, byte_we, byte_load, slt, lui, addm;
    input  [5:0] opcode, funct;
    input        zero;
    //from lab5
    wire inst_addi = opcode == `OP_ADDI;
    wire inst_andi = opcode == `OP_ANDI;
    wire inst_ori = opcode == `OP_ORI;
    wire inst_xori = opcode == `OP_XORI;
    wire inst_add = (opcode == `OP_OTHER0 ) & (funct == `OP0_ADD);
    wire inst_sub = (opcode == `OP_OTHER0 ) & (funct == `OP0_SUB);
    wire inst_and = (opcode == `OP_OTHER0 ) & (funct == `OP0_AND);
    wire inst_or  = (opcode == `OP_OTHER0 ) & (funct == `OP0_OR);
    wire inst_nor = (opcode == `OP_OTHER0 ) & (funct == `OP0_NOR);
    wire inst_xor = (opcode == `OP_OTHER0 ) & (funct == `OP0_XOR);
    //lab6 new
    wire inst_beq = (opcode == `OP_BEQ) & (zero == 1);
    wire inst_bne = (opcode == `OP_BNE) & (zero == 0);
    wire inst_beq_bne_false = ((opcode == `OP_BEQ)/* & (zero == 0)*/) | ((opcode == `OP_BNE)/* & (zero == 1)*/);
    wire inst_j = opcode == `OP_J;
    wire inst_jr = (opcode == `OP_OTHER0 ) & (funct == `OP0_JR);
    wire inst_lui = opcode == `OP_LUI;
    wire inst_slt = (opcode == `OP_OTHER0 ) & (funct == `OP0_SLT);
    wire inst_lw = opcode == `OP_LW;
    wire inst_lbu = opcode == `OP_LBU;
    wire inst_sw = opcode == `OP_SW;
    wire inst_sb = opcode == `OP_SB;
    wire inst_addm = (opcode == `OP_OTHER0 ) & (funct == `OP0_ADDM);

    //assigning all don't cares to 0
    assign alu_op = inst_add ? 3'b010 :
    inst_sub ? 3'b011 :
    inst_and ? 3'b100 :
    inst_or ? 3'b101 :
    inst_nor ? 3'b110 :
    inst_xor ? 3'b111 :
    inst_addi ? 3'b010 :
    inst_andi ? 3'b100 :
    inst_ori ? 3'b101 :
    inst_xori ? 3'b111:

    inst_beq ? 3'b011:
    inst_bne ? 3'b011:
    inst_beq_bne_false ? 3'b011:
    inst_slt ? 3'b011:
    inst_lw ? 3'b010:
    inst_lbu ? 3'b010:
    inst_sw ? 3'b010:
    inst_sb ? 3'b010:
    inst_addm ? 3'b010:
    3'b000;

    assign rd_src =
    inst_addi ? 1 :
    inst_andi ? 1 :
    inst_ori ? 1 :
    inst_xori ? 1:

    inst_beq ? 1:
    inst_bne ? 1:
    inst_lui ? 1:
    inst_lw ? 1:
    inst_lbu ? 1:
    inst_sw ? 1:
    inst_sb ? 1:
    0;

    assign alu_src2 =
    inst_addi ? 1 :
    inst_andi ? 1 :
    inst_ori ? 1 :
    inst_xori ? 1:

    inst_lw ? 1 :
    inst_lbu ? 1 :
    inst_sw ? 1 :
    inst_sb ? 1:
    0;


    assign writeenable = inst_add | inst_sub | inst_and |inst_or |inst_nor| inst_xor | inst_addi |inst_andi|inst_ori|inst_xori
                    | inst_lui | inst_slt | inst_lw | inst_lbu | inst_addm;
    assign except = ~writeenable & ~inst_beq & ~inst_bne & ~inst_beq_bne_false & ~inst_j & ~inst_jr & ~inst_sw & ~inst_sb;

    assign control_type[0] = inst_beq ? 1 :
    inst_bne ? 1 :
    inst_jr ? 1 :
    0;
    assign control_type[1] = inst_j ? 1 :
    inst_jr ? 1 :
    0;

    assign mem_read = inst_lw | inst_lbu;
    assign word_we = inst_sw;
    assign byte_we = inst_sb;
    assign byte_load = inst_lbu;
    assign lui = inst_lui;
    assign slt = inst_slt;
    assign addm = inst_addm;

endmodule // mips_decode
